// pd_block.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module pd_block (
		input  wire        clock_clk,                //            clock.clk
		input  wire        clock_sreset_reset_n,     //     clock_sreset.reset_n
		output wire [9:0]  led_export,               //              led.export
		output wire [12:0] sdram_addr,               //            sdram.addr
		output wire [1:0]  sdram_ba,                 //                 .ba
		output wire        sdram_cas_n,              //                 .cas_n
		output wire        sdram_cke,                //                 .cke
		output wire        sdram_cs_n,               //                 .cs_n
		inout  wire [15:0] sdram_dq,                 //                 .dq
		output wire [1:0]  sdram_dqm,                //                 .dqm
		output wire        sdram_ras_n,              //                 .ras_n
		output wire        sdram_we_n,               //                 .we_n
		output wire [15:0] vga_rgb,                  //              vga.rgb
		output wire        vga_valid,                //                 .valid
		output wire        vga_vsync,                //                 .vsync
		output wire        vga_hsync,                //                 .hsync
		input  wire        vga_clock_clk,            //        vga_clock.clk
		input  wire        vga_clock_sreset_reset_n  // vga_clock_sreset.reset_n
	);

	wire         frame_reader_source_valid;                                 // frame_reader:st_valid -> vga_out:st_valid
	wire  [15:0] frame_reader_source_data;                                  // frame_reader:st_data -> vga_out:st_data
	wire         frame_reader_source_ready;                                 // vga_out:st_ready -> frame_reader:st_ready
	wire         frame_reader_source_startofpacket;                         // frame_reader:st_sop -> vga_out:st_sop
	wire         frame_reader_source_endofpacket;                           // frame_reader:st_eop -> vga_out:st_eop
	wire         from_memory1_source_valid;                                 // from_memory1:st_valid -> pad1:si_valid
	wire  [15:0] from_memory1_source_data;                                  // from_memory1:st_data -> pad1:si_data
	wire         from_memory1_source_ready;                                 // pad1:si_ready -> from_memory1:st_ready
	wire         from_memory1_source_startofpacket;                         // from_memory1:st_sop -> pad1:si_sop
	wire         from_memory1_source_endofpacket;                           // from_memory1:st_eop -> pad1:si_eop
	wire         pad1_source_valid;                                         // pad1:so_valid -> conv1:st_valid
	wire  [15:0] pad1_source_data;                                          // pad1:so_data -> conv1:st_data
	wire         pad1_source_ready;                                         // conv1:st_ready -> pad1:so_ready
	wire         pad1_source_startofpacket;                                 // pad1:so_sop -> conv1:st_sop
	wire         pad1_source_endofpacket;                                   // pad1:so_eop -> conv1:st_eop
	wire  [15:0] rgb_tensor_avalon_master_readdata;                         // mm_interconnect_0:rgb_tensor_avalon_master_readdata -> rgb_tensor:m_readdata
	wire         rgb_tensor_avalon_master_waitrequest;                      // mm_interconnect_0:rgb_tensor_avalon_master_waitrequest -> rgb_tensor:m_waitrequest
	wire  [31:0] rgb_tensor_avalon_master_address;                          // rgb_tensor:m_address -> mm_interconnect_0:rgb_tensor_avalon_master_address
	wire   [1:0] rgb_tensor_avalon_master_byteenable;                       // rgb_tensor:m_byteenable -> mm_interconnect_0:rgb_tensor_avalon_master_byteenable
	wire         rgb_tensor_avalon_master_read;                             // rgb_tensor:m_read -> mm_interconnect_0:rgb_tensor_avalon_master_read
	wire  [15:0] rgb_tensor_avalon_master_writedata;                        // rgb_tensor:m_writedata -> mm_interconnect_0:rgb_tensor_avalon_master_writedata
	wire         rgb_tensor_avalon_master_write;                            // rgb_tensor:m_write -> mm_interconnect_0:rgb_tensor_avalon_master_write
	wire  [31:0] nios2e_data_master_readdata;                               // mm_interconnect_0:nios2e_data_master_readdata -> nios2e:d_readdata
	wire         nios2e_data_master_waitrequest;                            // mm_interconnect_0:nios2e_data_master_waitrequest -> nios2e:d_waitrequest
	wire         nios2e_data_master_debugaccess;                            // nios2e:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2e_data_master_debugaccess
	wire  [27:0] nios2e_data_master_address;                                // nios2e:d_address -> mm_interconnect_0:nios2e_data_master_address
	wire   [3:0] nios2e_data_master_byteenable;                             // nios2e:d_byteenable -> mm_interconnect_0:nios2e_data_master_byteenable
	wire         nios2e_data_master_read;                                   // nios2e:d_read -> mm_interconnect_0:nios2e_data_master_read
	wire         nios2e_data_master_write;                                  // nios2e:d_write -> mm_interconnect_0:nios2e_data_master_write
	wire  [31:0] nios2e_data_master_writedata;                              // nios2e:d_writedata -> mm_interconnect_0:nios2e_data_master_writedata
	wire  [31:0] nios2e_instruction_master_readdata;                        // mm_interconnect_0:nios2e_instruction_master_readdata -> nios2e:i_readdata
	wire         nios2e_instruction_master_waitrequest;                     // mm_interconnect_0:nios2e_instruction_master_waitrequest -> nios2e:i_waitrequest
	wire  [27:0] nios2e_instruction_master_address;                         // nios2e:i_address -> mm_interconnect_0:nios2e_instruction_master_address
	wire         nios2e_instruction_master_read;                            // nios2e:i_read -> mm_interconnect_0:nios2e_instruction_master_read
	wire  [15:0] from_memory1_read_master_readdata;                         // mm_interconnect_0:from_memory1_read_master_readdata -> from_memory1:rm_readdata
	wire         from_memory1_read_master_waitrequest;                      // mm_interconnect_0:from_memory1_read_master_waitrequest -> from_memory1:rm_waitrequest
	wire  [31:0] from_memory1_read_master_address;                          // from_memory1:rm_address -> mm_interconnect_0:from_memory1_read_master_address
	wire   [1:0] from_memory1_read_master_byteenable;                       // from_memory1:rm_byteenable -> mm_interconnect_0:from_memory1_read_master_byteenable
	wire         from_memory1_read_master_read;                             // from_memory1:rm_read -> mm_interconnect_0:from_memory1_read_master_read
	wire         from_memory1_read_master_readdatavalid;                    // mm_interconnect_0:from_memory1_read_master_readdatavalid -> from_memory1:rm_readdatavalid
	wire  [15:0] dma_read_master_readdata;                                  // mm_interconnect_0:dma_read_master_readdata -> dma:mr_readdata
	wire         dma_read_master_waitrequest;                               // mm_interconnect_0:dma_read_master_waitrequest -> dma:mr_waitrequest
	wire  [31:0] dma_read_master_address;                                   // dma:mr_address -> mm_interconnect_0:dma_read_master_address
	wire   [1:0] dma_read_master_byteenable;                                // dma:mr_byteenable -> mm_interconnect_0:dma_read_master_byteenable
	wire         dma_read_master_read;                                      // dma:mr_read -> mm_interconnect_0:dma_read_master_read
	wire         dma_write_master_waitrequest;                              // mm_interconnect_0:dma_write_master_waitrequest -> dma:mw_waitrequest
	wire  [31:0] dma_write_master_address;                                  // dma:mw_address -> mm_interconnect_0:dma_write_master_address
	wire   [1:0] dma_write_master_byteenable;                               // dma:mw_byteenable -> mm_interconnect_0:dma_write_master_byteenable
	wire         dma_write_master_write;                                    // dma:mw_write -> mm_interconnect_0:dma_write_master_write
	wire  [15:0] dma_write_master_writedata;                                // dma:mw_writedata -> mm_interconnect_0:dma_write_master_writedata
	wire  [15:0] mm_interconnect_0_bridge2_s0_readdata;                     // bridge2:s0_readdata -> mm_interconnect_0:bridge2_s0_readdata
	wire         mm_interconnect_0_bridge2_s0_waitrequest;                  // bridge2:s0_waitrequest -> mm_interconnect_0:bridge2_s0_waitrequest
	wire         mm_interconnect_0_bridge2_s0_debugaccess;                  // mm_interconnect_0:bridge2_s0_debugaccess -> bridge2:s0_debugaccess
	wire  [26:0] mm_interconnect_0_bridge2_s0_address;                      // mm_interconnect_0:bridge2_s0_address -> bridge2:s0_address
	wire         mm_interconnect_0_bridge2_s0_read;                         // mm_interconnect_0:bridge2_s0_read -> bridge2:s0_read
	wire   [1:0] mm_interconnect_0_bridge2_s0_byteenable;                   // mm_interconnect_0:bridge2_s0_byteenable -> bridge2:s0_byteenable
	wire         mm_interconnect_0_bridge2_s0_readdatavalid;                // bridge2:s0_readdatavalid -> mm_interconnect_0:bridge2_s0_readdatavalid
	wire         mm_interconnect_0_bridge2_s0_write;                        // mm_interconnect_0:bridge2_s0_write -> bridge2:s0_write
	wire  [15:0] mm_interconnect_0_bridge2_s0_writedata;                    // mm_interconnect_0:bridge2_s0_writedata -> bridge2:s0_writedata
	wire   [5:0] mm_interconnect_0_bridge2_s0_burstcount;                   // mm_interconnect_0:bridge2_s0_burstcount -> bridge2:s0_burstcount
	wire  [31:0] mm_interconnect_0_nios2e_debug_mem_slave_readdata;         // nios2e:debug_mem_slave_readdata -> mm_interconnect_0:nios2e_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2e_debug_mem_slave_waitrequest;      // nios2e:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2e_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2e_debug_mem_slave_debugaccess;      // mm_interconnect_0:nios2e_debug_mem_slave_debugaccess -> nios2e:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2e_debug_mem_slave_address;          // mm_interconnect_0:nios2e_debug_mem_slave_address -> nios2e:debug_mem_slave_address
	wire         mm_interconnect_0_nios2e_debug_mem_slave_read;             // mm_interconnect_0:nios2e_debug_mem_slave_read -> nios2e:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2e_debug_mem_slave_byteenable;       // mm_interconnect_0:nios2e_debug_mem_slave_byteenable -> nios2e:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2e_debug_mem_slave_write;            // mm_interconnect_0:nios2e_debug_mem_slave_write -> nios2e:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2e_debug_mem_slave_writedata;        // mm_interconnect_0:nios2e_debug_mem_slave_writedata -> nios2e:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_ram_s1_chipselect;                // mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_readdata;                  // onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	wire  [11:0] mm_interconnect_0_onchip_ram_s1_address;                   // mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	wire   [3:0] mm_interconnect_0_onchip_ram_s1_byteenable;                // mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	wire         mm_interconnect_0_onchip_ram_s1_write;                     // mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_writedata;                 // mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	wire         mm_interconnect_0_onchip_ram_s1_clken;                     // mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_bridge1_s0_readdata;                     // bridge1:s0_readdata -> mm_interconnect_0:bridge1_s0_readdata
	wire         mm_interconnect_0_bridge1_s0_waitrequest;                  // bridge1:s0_waitrequest -> mm_interconnect_0:bridge1_s0_waitrequest
	wire         mm_interconnect_0_bridge1_s0_debugaccess;                  // mm_interconnect_0:bridge1_s0_debugaccess -> bridge1:s0_debugaccess
	wire   [7:0] mm_interconnect_0_bridge1_s0_address;                      // mm_interconnect_0:bridge1_s0_address -> bridge1:s0_address
	wire         mm_interconnect_0_bridge1_s0_read;                         // mm_interconnect_0:bridge1_s0_read -> bridge1:s0_read
	wire   [3:0] mm_interconnect_0_bridge1_s0_byteenable;                   // mm_interconnect_0:bridge1_s0_byteenable -> bridge1:s0_byteenable
	wire         mm_interconnect_0_bridge1_s0_readdatavalid;                // bridge1:s0_readdatavalid -> mm_interconnect_0:bridge1_s0_readdatavalid
	wire         mm_interconnect_0_bridge1_s0_write;                        // mm_interconnect_0:bridge1_s0_write -> bridge1:s0_write
	wire  [31:0] mm_interconnect_0_bridge1_s0_writedata;                    // mm_interconnect_0:bridge1_s0_writedata -> bridge1:s0_writedata
	wire   [4:0] mm_interconnect_0_bridge1_s0_burstcount;                   // mm_interconnect_0:bridge1_s0_burstcount -> bridge1:s0_burstcount
	wire         mm_interconnect_0_led_s1_chipselect;                       // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                         // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;                          // mm_interconnect_0:led_s1_address -> led:address
	wire         mm_interconnect_0_led_s1_write;                            // mm_interconnect_0:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                        // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire  [31:0] mm_interconnect_0_frame_reader_slave_readdata;             // frame_reader:s_readdata -> mm_interconnect_0:frame_reader_slave_readdata
	wire         mm_interconnect_0_frame_reader_slave_waitrequest;          // frame_reader:s_waitrequest -> mm_interconnect_0:frame_reader_slave_waitrequest
	wire   [3:0] mm_interconnect_0_frame_reader_slave_address;              // mm_interconnect_0:frame_reader_slave_address -> frame_reader:s_address
	wire         mm_interconnect_0_frame_reader_slave_read;                 // mm_interconnect_0:frame_reader_slave_read -> frame_reader:s_read
	wire         mm_interconnect_0_frame_reader_slave_write;                // mm_interconnect_0:frame_reader_slave_write -> frame_reader:s_write
	wire  [31:0] mm_interconnect_0_frame_reader_slave_writedata;            // mm_interconnect_0:frame_reader_slave_writedata -> frame_reader:s_writedata
	wire  [31:0] mm_interconnect_0_vga_out_slave_readdata;                  // vga_out:s_readdata -> mm_interconnect_0:vga_out_slave_readdata
	wire         mm_interconnect_0_vga_out_slave_waitrequest;               // vga_out:s_waitrequest -> mm_interconnect_0:vga_out_slave_waitrequest
	wire   [3:0] mm_interconnect_0_vga_out_slave_address;                   // mm_interconnect_0:vga_out_slave_address -> vga_out:s_address
	wire         mm_interconnect_0_vga_out_slave_read;                      // mm_interconnect_0:vga_out_slave_read -> vga_out:s_read
	wire         mm_interconnect_0_vga_out_slave_write;                     // mm_interconnect_0:vga_out_slave_write -> vga_out:s_write
	wire  [31:0] mm_interconnect_0_vga_out_slave_writedata;                 // mm_interconnect_0:vga_out_slave_writedata -> vga_out:s_writedata
	wire         bridge2_m0_waitrequest;                                    // mm_interconnect_1:bridge2_m0_waitrequest -> bridge2:m0_waitrequest
	wire  [15:0] bridge2_m0_readdata;                                       // mm_interconnect_1:bridge2_m0_readdata -> bridge2:m0_readdata
	wire         bridge2_m0_debugaccess;                                    // bridge2:m0_debugaccess -> mm_interconnect_1:bridge2_m0_debugaccess
	wire  [26:0] bridge2_m0_address;                                        // bridge2:m0_address -> mm_interconnect_1:bridge2_m0_address
	wire         bridge2_m0_read;                                           // bridge2:m0_read -> mm_interconnect_1:bridge2_m0_read
	wire   [1:0] bridge2_m0_byteenable;                                     // bridge2:m0_byteenable -> mm_interconnect_1:bridge2_m0_byteenable
	wire         bridge2_m0_readdatavalid;                                  // mm_interconnect_1:bridge2_m0_readdatavalid -> bridge2:m0_readdatavalid
	wire  [15:0] bridge2_m0_writedata;                                      // bridge2:m0_writedata -> mm_interconnect_1:bridge2_m0_writedata
	wire         bridge2_m0_write;                                          // bridge2:m0_write -> mm_interconnect_1:bridge2_m0_write
	wire   [5:0] bridge2_m0_burstcount;                                     // bridge2:m0_burstcount -> mm_interconnect_1:bridge2_m0_burstcount
	wire  [15:0] frame_reader_read_master_readdata;                         // mm_interconnect_1:frame_reader_read_master_readdata -> frame_reader:m_readdata
	wire         frame_reader_read_master_waitrequest;                      // mm_interconnect_1:frame_reader_read_master_waitrequest -> frame_reader:m_waitrequest
	wire  [31:0] frame_reader_read_master_address;                          // frame_reader:m_address -> mm_interconnect_1:frame_reader_read_master_address
	wire   [1:0] frame_reader_read_master_byteenable;                       // frame_reader:m_byteenable -> mm_interconnect_1:frame_reader_read_master_byteenable
	wire         frame_reader_read_master_read;                             // frame_reader:m_read -> mm_interconnect_1:frame_reader_read_master_read
	wire         frame_reader_read_master_readdatavalid;                    // mm_interconnect_1:frame_reader_read_master_readdatavalid -> frame_reader:m_readdatavalid
	wire         mm_interconnect_1_sdram_s1_chipselect;                     // mm_interconnect_1:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_1_sdram_s1_readdata;                       // sdram:za_data -> mm_interconnect_1:sdram_s1_readdata
	wire         mm_interconnect_1_sdram_s1_waitrequest;                    // sdram:za_waitrequest -> mm_interconnect_1:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_1_sdram_s1_address;                        // mm_interconnect_1:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_1_sdram_s1_read;                           // mm_interconnect_1:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_1_sdram_s1_byteenable;                     // mm_interconnect_1:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_1_sdram_s1_readdatavalid;                  // sdram:za_valid -> mm_interconnect_1:sdram_s1_readdatavalid
	wire         mm_interconnect_1_sdram_s1_write;                          // mm_interconnect_1:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_1_sdram_s1_writedata;                      // mm_interconnect_1:sdram_s1_writedata -> sdram:az_data
	wire         bridge1_m0_waitrequest;                                    // mm_interconnect_2:bridge1_m0_waitrequest -> bridge1:m0_waitrequest
	wire  [31:0] bridge1_m0_readdata;                                       // mm_interconnect_2:bridge1_m0_readdata -> bridge1:m0_readdata
	wire         bridge1_m0_debugaccess;                                    // bridge1:m0_debugaccess -> mm_interconnect_2:bridge1_m0_debugaccess
	wire   [7:0] bridge1_m0_address;                                        // bridge1:m0_address -> mm_interconnect_2:bridge1_m0_address
	wire         bridge1_m0_read;                                           // bridge1:m0_read -> mm_interconnect_2:bridge1_m0_read
	wire   [3:0] bridge1_m0_byteenable;                                     // bridge1:m0_byteenable -> mm_interconnect_2:bridge1_m0_byteenable
	wire         bridge1_m0_readdatavalid;                                  // mm_interconnect_2:bridge1_m0_readdatavalid -> bridge1:m0_readdatavalid
	wire  [31:0] bridge1_m0_writedata;                                      // bridge1:m0_writedata -> mm_interconnect_2:bridge1_m0_writedata
	wire         bridge1_m0_write;                                          // bridge1:m0_write -> mm_interconnect_2:bridge1_m0_write
	wire   [4:0] bridge1_m0_burstcount;                                     // bridge1:m0_burstcount -> mm_interconnect_2:bridge1_m0_burstcount
	wire  [31:0] mm_interconnect_2_dma_slave_readdata;                      // dma:s_readdata -> mm_interconnect_2:dma_slave_readdata
	wire         mm_interconnect_2_dma_slave_waitrequest;                   // dma:s_waitrequest -> mm_interconnect_2:dma_slave_waitrequest
	wire   [3:0] mm_interconnect_2_dma_slave_address;                       // mm_interconnect_2:dma_slave_address -> dma:s_address
	wire         mm_interconnect_2_dma_slave_read;                          // mm_interconnect_2:dma_slave_read -> dma:s_read
	wire         mm_interconnect_2_dma_slave_write;                         // mm_interconnect_2:dma_slave_write -> dma:s_write
	wire  [31:0] mm_interconnect_2_dma_slave_writedata;                     // mm_interconnect_2:dma_slave_writedata -> dma:s_writedata
	wire  [31:0] mm_interconnect_2_rgb_tensor_slave_readdata;               // rgb_tensor:s_readdata -> mm_interconnect_2:rgb_tensor_slave_readdata
	wire         mm_interconnect_2_rgb_tensor_slave_waitrequest;            // rgb_tensor:s_waitrequest -> mm_interconnect_2:rgb_tensor_slave_waitrequest
	wire   [3:0] mm_interconnect_2_rgb_tensor_slave_address;                // mm_interconnect_2:rgb_tensor_slave_address -> rgb_tensor:s_address
	wire         mm_interconnect_2_rgb_tensor_slave_read;                   // mm_interconnect_2:rgb_tensor_slave_read -> rgb_tensor:s_read
	wire         mm_interconnect_2_rgb_tensor_slave_write;                  // mm_interconnect_2:rgb_tensor_slave_write -> rgb_tensor:s_write
	wire  [31:0] mm_interconnect_2_rgb_tensor_slave_writedata;              // mm_interconnect_2:rgb_tensor_slave_writedata -> rgb_tensor:s_writedata
	wire  [31:0] mm_interconnect_2_from_memory1_slave_readdata;             // from_memory1:s_readdata -> mm_interconnect_2:from_memory1_slave_readdata
	wire         mm_interconnect_2_from_memory1_slave_waitrequest;          // from_memory1:s_waitrequest -> mm_interconnect_2:from_memory1_slave_waitrequest
	wire   [3:0] mm_interconnect_2_from_memory1_slave_address;              // mm_interconnect_2:from_memory1_slave_address -> from_memory1:s_address
	wire         mm_interconnect_2_from_memory1_slave_read;                 // mm_interconnect_2:from_memory1_slave_read -> from_memory1:s_read
	wire         mm_interconnect_2_from_memory1_slave_write;                // mm_interconnect_2:from_memory1_slave_write -> from_memory1:s_write
	wire  [31:0] mm_interconnect_2_from_memory1_slave_writedata;            // mm_interconnect_2:from_memory1_slave_writedata -> from_memory1:s_writedata
	wire         mm_interconnect_2_conv1_slave_waitrequest;                 // conv1:s_waitrequest -> mm_interconnect_2:conv1_slave_waitrequest
	wire   [0:0] mm_interconnect_2_conv1_slave_address;                     // mm_interconnect_2:conv1_slave_address -> conv1:s_address
	wire         mm_interconnect_2_conv1_slave_write;                       // mm_interconnect_2:conv1_slave_write -> conv1:s_write
	wire  [15:0] mm_interconnect_2_conv1_slave_writedata;                   // mm_interconnect_2:conv1_slave_writedata -> conv1:s_writedata
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // dma:s_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2e_irq_irq;                                            // irq_mapper:sender_irq -> nios2e:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [bridge1:reset, bridge2:reset, conv1:clock_sreset, from_memory1:clock_sreset, irq_mapper:reset, jtag_uart:rst_n, led:reset_n, mm_interconnect_0:nios2e_reset_reset_bridge_in_reset_reset, mm_interconnect_0:rgb_tensor_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:bridge2_reset_reset_bridge_in_reset_reset, mm_interconnect_1:frame_reader_clock_sreset_reset_bridge_in_reset_reset, mm_interconnect_2:bridge1_reset_reset_bridge_in_reset_reset, mm_interconnect_2:rgb_tensor_reset_sink_reset_bridge_in_reset_reset, nios2e:reset_n, onchip_ram:reset, pad1:clock_sreset, rst_translator:in_reset, sdram:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [nios2e:reset_req, onchip_ram:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> dma:clock_sreset
	wire         nios2e_debug_reset_request_reset;                          // nios2e:debug_reset_request -> [rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_002_reset_out_reset;                        // rst_controller_002:reset_out -> [mm_interconnect_0:dma_clock_sreset_reset_bridge_in_reset_reset, mm_interconnect_0:dma_read_master_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_2:dma_clock_sreset_reset_bridge_in_reset_reset, mm_interconnect_2:dma_slave_translator_reset_reset_bridge_in_reset_reset]

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (8),
		.BURSTCOUNT_WIDTH  (5),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) bridge1 (
		.clk              (clock_clk),                                  //   clk.clk
		.reset            (rst_controller_reset_out_reset),             // reset.reset
		.s0_waitrequest   (mm_interconnect_0_bridge1_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_bridge1_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_bridge1_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_bridge1_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_bridge1_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_bridge1_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_bridge1_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_bridge1_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_bridge1_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_bridge1_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (bridge1_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (bridge1_m0_readdata),                        //      .readdata
		.m0_readdatavalid (bridge1_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (bridge1_m0_burstcount),                      //      .burstcount
		.m0_writedata     (bridge1_m0_writedata),                       //      .writedata
		.m0_address       (bridge1_m0_address),                         //      .address
		.m0_write         (bridge1_m0_write),                           //      .write
		.m0_read          (bridge1_m0_read),                            //      .read
		.m0_byteenable    (bridge1_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (bridge1_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                           // (terminated)
		.m0_response      (2'b00)                                       // (terminated)
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (16),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (27),
		.BURSTCOUNT_WIDTH  (6),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) bridge2 (
		.clk              (clock_clk),                                  //   clk.clk
		.reset            (rst_controller_reset_out_reset),             // reset.reset
		.s0_waitrequest   (mm_interconnect_0_bridge2_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_bridge2_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_bridge2_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_bridge2_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_bridge2_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_bridge2_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_bridge2_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_bridge2_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_bridge2_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_bridge2_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (bridge2_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (bridge2_m0_readdata),                        //      .readdata
		.m0_readdatavalid (bridge2_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (bridge2_m0_burstcount),                      //      .burstcount
		.m0_writedata     (bridge2_m0_writedata),                       //      .writedata
		.m0_address       (bridge2_m0_address),                         //      .address
		.m0_write         (bridge2_m0_write),                           //      .write
		.m0_read          (bridge2_m0_read),                            //      .read
		.m0_byteenable    (bridge2_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (bridge2_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                           // (terminated)
		.m0_response      (2'b00)                                       // (terminated)
	);

	convolution_calc #(
		.XRES        (64),
		.KX          (3),
		.KY          (3),
		.EXP         (8),
		.MANT        (7),
		.MLT_LCYCLES (1),
		.ADD_LCYCLES (4)
	) conv1 (
		.clock         (clock_clk),                                 //        clock.clk
		.clock_sreset  (rst_controller_reset_out_reset),            // clock_sreset.reset
		.result_valid  (),                                          //       source.valid
		.result        (),                                          //             .data
		.st_ready      (pad1_source_ready),                         //         sink.ready
		.st_valid      (pad1_source_valid),                         //             .valid
		.st_sop        (pad1_source_startofpacket),                 //             .startofpacket
		.st_eop        (pad1_source_endofpacket),                   //             .endofpacket
		.st_data       (pad1_source_data),                          //             .data
		.s_address     (mm_interconnect_2_conv1_slave_address),     //        slave.address
		.s_writedata   (mm_interconnect_2_conv1_slave_writedata),   //             .writedata
		.s_write       (mm_interconnect_2_conv1_slave_write),       //             .write
		.s_waitrequest (mm_interconnect_2_conv1_slave_waitrequest)  //             .waitrequest
	);

	dma_engine dma (
		.clock          (clock_clk),                               //        clock.clk
		.clock_sreset   (rst_controller_001_reset_out_reset),      // clock_sreset.reset
		.s_address      (mm_interconnect_2_dma_slave_address),     //        slave.address
		.s_writedata    (mm_interconnect_2_dma_slave_writedata),   //             .writedata
		.s_readdata     (mm_interconnect_2_dma_slave_readdata),    //             .readdata
		.s_read         (mm_interconnect_2_dma_slave_read),        //             .read
		.s_write        (mm_interconnect_2_dma_slave_write),       //             .write
		.s_waitrequest  (mm_interconnect_2_dma_slave_waitrequest), //             .waitrequest
		.s_irq          (irq_mapper_receiver1_irq),                //          irq.irq
		.mr_address     (dma_read_master_address),                 //  read_master.address
		.mr_byteenable  (dma_read_master_byteenable),              //             .byteenable
		.mr_readdata    (dma_read_master_readdata),                //             .readdata
		.mr_waitrequest (dma_read_master_waitrequest),             //             .waitrequest
		.mr_read        (dma_read_master_read),                    //             .read
		.mw_address     (dma_write_master_address),                // write_master.address
		.mw_byteenable  (dma_write_master_byteenable),             //             .byteenable
		.mw_write       (dma_write_master_write),                  //             .write
		.mw_writedata   (dma_write_master_writedata),              //             .writedata
		.mw_waitrequest (dma_write_master_waitrequest)             //             .waitrequest
	);

	frame_reader #(
		.XRES (640),
		.YRES (480)
	) frame_reader (
		.m_address       (frame_reader_read_master_address),                 //  read_master.address
		.m_byteenable    (frame_reader_read_master_byteenable),              //             .byteenable
		.m_readdata      (frame_reader_read_master_readdata),                //             .readdata
		.m_read          (frame_reader_read_master_read),                    //             .read
		.m_readdatavalid (frame_reader_read_master_readdatavalid),           //             .readdatavalid
		.m_waitrequest   (frame_reader_read_master_waitrequest),             //             .waitrequest
		.s_address       (mm_interconnect_0_frame_reader_slave_address),     //        slave.address
		.s_readdata      (mm_interconnect_0_frame_reader_slave_readdata),    //             .readdata
		.s_writedata     (mm_interconnect_0_frame_reader_slave_writedata),   //             .writedata
		.s_read          (mm_interconnect_0_frame_reader_slave_read),        //             .read
		.s_write         (mm_interconnect_0_frame_reader_slave_write),       //             .write
		.s_waitrequest   (mm_interconnect_0_frame_reader_slave_waitrequest), //             .waitrequest
		.st_ready        (frame_reader_source_ready),                        //       source.ready
		.st_valid        (frame_reader_source_valid),                        //             .valid
		.st_sop          (frame_reader_source_startofpacket),                //             .startofpacket
		.st_eop          (frame_reader_source_endofpacket),                  //             .endofpacket
		.st_data         (frame_reader_source_data),                         //             .data
		.clock           (clock_clk),                                        //        clock.clk
		.clock_sreset    (~clock_sreset_reset_n)                             // clock_sreset.reset
	);

	stream_from_memory from_memory1 (
		.clock            (clock_clk),                                        //        clock.clk
		.clock_sreset     (rst_controller_reset_out_reset),                   // clock_sreset.reset
		.st_ready         (from_memory1_source_ready),                        //       source.ready
		.st_valid         (from_memory1_source_valid),                        //             .valid
		.st_sop           (from_memory1_source_startofpacket),                //             .startofpacket
		.st_eop           (from_memory1_source_endofpacket),                  //             .endofpacket
		.st_data          (from_memory1_source_data),                         //             .data
		.s_address        (mm_interconnect_2_from_memory1_slave_address),     //        slave.address
		.s_readdata       (mm_interconnect_2_from_memory1_slave_readdata),    //             .readdata
		.s_writedata      (mm_interconnect_2_from_memory1_slave_writedata),   //             .writedata
		.s_read           (mm_interconnect_2_from_memory1_slave_read),        //             .read
		.s_write          (mm_interconnect_2_from_memory1_slave_write),       //             .write
		.s_waitrequest    (mm_interconnect_2_from_memory1_slave_waitrequest), //             .waitrequest
		.rm_address       (from_memory1_read_master_address),                 //  read_master.address
		.rm_readdata      (from_memory1_read_master_readdata),                //             .readdata
		.rm_byteenable    (from_memory1_read_master_byteenable),              //             .byteenable
		.rm_read          (from_memory1_read_master_read),                    //             .read
		.rm_waitrequest   (from_memory1_read_master_waitrequest),             //             .waitrequest
		.rm_readdatavalid (from_memory1_read_master_readdatavalid)            //             .readdatavalid
	);

	pd_block_jtag_uart jtag_uart (
		.clk            (clock_clk),                                                 //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	pd_block_led led (
		.clk        (clock_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                           // external_connection.export
	);

	pd_block_nios2e nios2e (
		.clk                                 (clock_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (nios2e_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2e_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2e_data_master_read),                              //                          .read
		.d_readdata                          (nios2e_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2e_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2e_data_master_write),                             //                          .write
		.d_writedata                         (nios2e_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2e_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2e_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2e_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2e_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2e_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2e_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2e_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2e_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2e_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2e_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2e_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2e_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2e_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2e_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2e_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                      // custom_instruction_master.readra
	);

	pd_block_onchip_ram onchip_ram (
		.clk        (clock_clk),                                  //   clk1.clk
		.address    (mm_interconnect_0_onchip_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                        // (terminated)
	);

	pad_stream #(
		.PAD (1)
	) pad1 (
		.clock        (clock_clk),                         //        clock.clk
		.clock_sreset (rst_controller_reset_out_reset),    // clock_sreset.reset
		.so_ready     (pad1_source_ready),                 //       source.ready
		.so_valid     (pad1_source_valid),                 //             .valid
		.so_sop       (pad1_source_startofpacket),         //             .startofpacket
		.so_eop       (pad1_source_endofpacket),           //             .endofpacket
		.so_data      (pad1_source_data),                  //             .data
		.si_ready     (from_memory1_source_ready),         //         sink.ready
		.si_valid     (from_memory1_source_valid),         //             .valid
		.si_sop       (from_memory1_source_startofpacket), //             .startofpacket
		.si_eop       (from_memory1_source_endofpacket),   //             .endofpacket
		.si_data      (from_memory1_source_data)           //             .data
	);

	rgb_to_tensor rgb_tensor (
		.s_address     (mm_interconnect_2_rgb_tensor_slave_address),     //         slave.address
		.s_readdata    (mm_interconnect_2_rgb_tensor_slave_readdata),    //              .readdata
		.s_writedata   (mm_interconnect_2_rgb_tensor_slave_writedata),   //              .writedata
		.s_read        (mm_interconnect_2_rgb_tensor_slave_read),        //              .read
		.s_write       (mm_interconnect_2_rgb_tensor_slave_write),       //              .write
		.s_waitrequest (mm_interconnect_2_rgb_tensor_slave_waitrequest), //              .waitrequest
		.m_address     (rgb_tensor_avalon_master_address),               // avalon_master.address
		.m_writedata   (rgb_tensor_avalon_master_writedata),             //              .writedata
		.m_readdata    (rgb_tensor_avalon_master_readdata),              //              .readdata
		.m_byteenable  (rgb_tensor_avalon_master_byteenable),            //              .byteenable
		.m_read        (rgb_tensor_avalon_master_read),                  //              .read
		.m_write       (rgb_tensor_avalon_master_write),                 //              .write
		.m_waitrequest (rgb_tensor_avalon_master_waitrequest),           //              .waitrequest
		.clock         (clock_clk),                                      //    clock_sink.clk
		.clock_sreset  (~clock_sreset_reset_n)                           //    reset_sink.reset
	);

	pd_block_sdram sdram (
		.clk            (clock_clk),                                //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_1_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_1_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_1_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_1_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_1_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_1_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_1_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_1_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_1_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	vga_output #(
		.WIDTH         (16),
		.FIFO_DEPTH    (1024),
		.VGA_XRES      (640),
		.VGA_HSYNC     (96),
		.VGA_HFPORCH   (16),
		.VGA_HBPORCH   (48),
		.VGA_YRES      (480),
		.VGA_VSYNC     (2),
		.VGA_VFPORCH   (10),
		.VGA_VBPORCH   (33),
		.NO_SIGNAL_RGB (18'b001111111100000000)
	) vga_out (
		.st_ready         (frame_reader_source_ready),                   //             sink.ready
		.st_valid         (frame_reader_source_valid),                   //                 .valid
		.st_sop           (frame_reader_source_startofpacket),           //                 .startofpacket
		.st_eop           (frame_reader_source_endofpacket),             //                 .endofpacket
		.st_data          (frame_reader_source_data),                    //                 .data
		.clock            (clock_clk),                                   //            clock.clk
		.vga_rgb          (vga_rgb),                                     //              vga.rgb
		.vga_valid        (vga_valid),                                   //                 .valid
		.vga_vsync        (vga_vsync),                                   //                 .vsync
		.vga_hsync        (vga_hsync),                                   //                 .hsync
		.clock_sreset     (~clock_sreset_reset_n),                       //     clock_sreset.reset
		.vga_clock        (vga_clock_clk),                               //        vga_clock.clk
		.vga_clock_sreset (~vga_clock_sreset_reset_n),                   // vga_clock_sreset.reset
		.s_address        (mm_interconnect_0_vga_out_slave_address),     //            slave.address
		.s_writedata      (mm_interconnect_0_vga_out_slave_writedata),   //                 .writedata
		.s_readdata       (mm_interconnect_0_vga_out_slave_readdata),    //                 .readdata
		.s_read           (mm_interconnect_0_vga_out_slave_read),        //                 .read
		.s_write          (mm_interconnect_0_vga_out_slave_write),       //                 .write
		.s_waitrequest    (mm_interconnect_0_vga_out_slave_waitrequest)  //                 .waitrequest
	);

	pd_block_mm_interconnect_0 mm_interconnect_0 (
		.clock_clk_clk                                                (clock_clk),                                                 //                                              clock_clk.clk
		.dma_clock_sreset_reset_bridge_in_reset_reset                 (rst_controller_002_reset_out_reset),                        //                 dma_clock_sreset_reset_bridge_in_reset.reset
		.dma_read_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                        // dma_read_master_translator_reset_reset_bridge_in_reset.reset
		.nios2e_reset_reset_bridge_in_reset_reset                     (rst_controller_reset_out_reset),                            //                     nios2e_reset_reset_bridge_in_reset.reset
		.rgb_tensor_reset_sink_reset_bridge_in_reset_reset            (rst_controller_reset_out_reset),                            //            rgb_tensor_reset_sink_reset_bridge_in_reset.reset
		.dma_read_master_address                                      (dma_read_master_address),                                   //                                        dma_read_master.address
		.dma_read_master_waitrequest                                  (dma_read_master_waitrequest),                               //                                                       .waitrequest
		.dma_read_master_byteenable                                   (dma_read_master_byteenable),                                //                                                       .byteenable
		.dma_read_master_read                                         (dma_read_master_read),                                      //                                                       .read
		.dma_read_master_readdata                                     (dma_read_master_readdata),                                  //                                                       .readdata
		.dma_write_master_address                                     (dma_write_master_address),                                  //                                       dma_write_master.address
		.dma_write_master_waitrequest                                 (dma_write_master_waitrequest),                              //                                                       .waitrequest
		.dma_write_master_byteenable                                  (dma_write_master_byteenable),                               //                                                       .byteenable
		.dma_write_master_write                                       (dma_write_master_write),                                    //                                                       .write
		.dma_write_master_writedata                                   (dma_write_master_writedata),                                //                                                       .writedata
		.from_memory1_read_master_address                             (from_memory1_read_master_address),                          //                               from_memory1_read_master.address
		.from_memory1_read_master_waitrequest                         (from_memory1_read_master_waitrequest),                      //                                                       .waitrequest
		.from_memory1_read_master_byteenable                          (from_memory1_read_master_byteenable),                       //                                                       .byteenable
		.from_memory1_read_master_read                                (from_memory1_read_master_read),                             //                                                       .read
		.from_memory1_read_master_readdata                            (from_memory1_read_master_readdata),                         //                                                       .readdata
		.from_memory1_read_master_readdatavalid                       (from_memory1_read_master_readdatavalid),                    //                                                       .readdatavalid
		.nios2e_data_master_address                                   (nios2e_data_master_address),                                //                                     nios2e_data_master.address
		.nios2e_data_master_waitrequest                               (nios2e_data_master_waitrequest),                            //                                                       .waitrequest
		.nios2e_data_master_byteenable                                (nios2e_data_master_byteenable),                             //                                                       .byteenable
		.nios2e_data_master_read                                      (nios2e_data_master_read),                                   //                                                       .read
		.nios2e_data_master_readdata                                  (nios2e_data_master_readdata),                               //                                                       .readdata
		.nios2e_data_master_write                                     (nios2e_data_master_write),                                  //                                                       .write
		.nios2e_data_master_writedata                                 (nios2e_data_master_writedata),                              //                                                       .writedata
		.nios2e_data_master_debugaccess                               (nios2e_data_master_debugaccess),                            //                                                       .debugaccess
		.nios2e_instruction_master_address                            (nios2e_instruction_master_address),                         //                              nios2e_instruction_master.address
		.nios2e_instruction_master_waitrequest                        (nios2e_instruction_master_waitrequest),                     //                                                       .waitrequest
		.nios2e_instruction_master_read                               (nios2e_instruction_master_read),                            //                                                       .read
		.nios2e_instruction_master_readdata                           (nios2e_instruction_master_readdata),                        //                                                       .readdata
		.rgb_tensor_avalon_master_address                             (rgb_tensor_avalon_master_address),                          //                               rgb_tensor_avalon_master.address
		.rgb_tensor_avalon_master_waitrequest                         (rgb_tensor_avalon_master_waitrequest),                      //                                                       .waitrequest
		.rgb_tensor_avalon_master_byteenable                          (rgb_tensor_avalon_master_byteenable),                       //                                                       .byteenable
		.rgb_tensor_avalon_master_read                                (rgb_tensor_avalon_master_read),                             //                                                       .read
		.rgb_tensor_avalon_master_readdata                            (rgb_tensor_avalon_master_readdata),                         //                                                       .readdata
		.rgb_tensor_avalon_master_write                               (rgb_tensor_avalon_master_write),                            //                                                       .write
		.rgb_tensor_avalon_master_writedata                           (rgb_tensor_avalon_master_writedata),                        //                                                       .writedata
		.bridge1_s0_address                                           (mm_interconnect_0_bridge1_s0_address),                      //                                             bridge1_s0.address
		.bridge1_s0_write                                             (mm_interconnect_0_bridge1_s0_write),                        //                                                       .write
		.bridge1_s0_read                                              (mm_interconnect_0_bridge1_s0_read),                         //                                                       .read
		.bridge1_s0_readdata                                          (mm_interconnect_0_bridge1_s0_readdata),                     //                                                       .readdata
		.bridge1_s0_writedata                                         (mm_interconnect_0_bridge1_s0_writedata),                    //                                                       .writedata
		.bridge1_s0_burstcount                                        (mm_interconnect_0_bridge1_s0_burstcount),                   //                                                       .burstcount
		.bridge1_s0_byteenable                                        (mm_interconnect_0_bridge1_s0_byteenable),                   //                                                       .byteenable
		.bridge1_s0_readdatavalid                                     (mm_interconnect_0_bridge1_s0_readdatavalid),                //                                                       .readdatavalid
		.bridge1_s0_waitrequest                                       (mm_interconnect_0_bridge1_s0_waitrequest),                  //                                                       .waitrequest
		.bridge1_s0_debugaccess                                       (mm_interconnect_0_bridge1_s0_debugaccess),                  //                                                       .debugaccess
		.bridge2_s0_address                                           (mm_interconnect_0_bridge2_s0_address),                      //                                             bridge2_s0.address
		.bridge2_s0_write                                             (mm_interconnect_0_bridge2_s0_write),                        //                                                       .write
		.bridge2_s0_read                                              (mm_interconnect_0_bridge2_s0_read),                         //                                                       .read
		.bridge2_s0_readdata                                          (mm_interconnect_0_bridge2_s0_readdata),                     //                                                       .readdata
		.bridge2_s0_writedata                                         (mm_interconnect_0_bridge2_s0_writedata),                    //                                                       .writedata
		.bridge2_s0_burstcount                                        (mm_interconnect_0_bridge2_s0_burstcount),                   //                                                       .burstcount
		.bridge2_s0_byteenable                                        (mm_interconnect_0_bridge2_s0_byteenable),                   //                                                       .byteenable
		.bridge2_s0_readdatavalid                                     (mm_interconnect_0_bridge2_s0_readdatavalid),                //                                                       .readdatavalid
		.bridge2_s0_waitrequest                                       (mm_interconnect_0_bridge2_s0_waitrequest),                  //                                                       .waitrequest
		.bridge2_s0_debugaccess                                       (mm_interconnect_0_bridge2_s0_debugaccess),                  //                                                       .debugaccess
		.frame_reader_slave_address                                   (mm_interconnect_0_frame_reader_slave_address),              //                                     frame_reader_slave.address
		.frame_reader_slave_write                                     (mm_interconnect_0_frame_reader_slave_write),                //                                                       .write
		.frame_reader_slave_read                                      (mm_interconnect_0_frame_reader_slave_read),                 //                                                       .read
		.frame_reader_slave_readdata                                  (mm_interconnect_0_frame_reader_slave_readdata),             //                                                       .readdata
		.frame_reader_slave_writedata                                 (mm_interconnect_0_frame_reader_slave_writedata),            //                                                       .writedata
		.frame_reader_slave_waitrequest                               (mm_interconnect_0_frame_reader_slave_waitrequest),          //                                                       .waitrequest
		.jtag_uart_avalon_jtag_slave_address                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                            jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                                       .write
		.jtag_uart_avalon_jtag_slave_read                             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                                       .read
		.jtag_uart_avalon_jtag_slave_readdata                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                                       .readdata
		.jtag_uart_avalon_jtag_slave_writedata                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                                       .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                                       .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                                       .chipselect
		.led_s1_address                                               (mm_interconnect_0_led_s1_address),                          //                                                 led_s1.address
		.led_s1_write                                                 (mm_interconnect_0_led_s1_write),                            //                                                       .write
		.led_s1_readdata                                              (mm_interconnect_0_led_s1_readdata),                         //                                                       .readdata
		.led_s1_writedata                                             (mm_interconnect_0_led_s1_writedata),                        //                                                       .writedata
		.led_s1_chipselect                                            (mm_interconnect_0_led_s1_chipselect),                       //                                                       .chipselect
		.nios2e_debug_mem_slave_address                               (mm_interconnect_0_nios2e_debug_mem_slave_address),          //                                 nios2e_debug_mem_slave.address
		.nios2e_debug_mem_slave_write                                 (mm_interconnect_0_nios2e_debug_mem_slave_write),            //                                                       .write
		.nios2e_debug_mem_slave_read                                  (mm_interconnect_0_nios2e_debug_mem_slave_read),             //                                                       .read
		.nios2e_debug_mem_slave_readdata                              (mm_interconnect_0_nios2e_debug_mem_slave_readdata),         //                                                       .readdata
		.nios2e_debug_mem_slave_writedata                             (mm_interconnect_0_nios2e_debug_mem_slave_writedata),        //                                                       .writedata
		.nios2e_debug_mem_slave_byteenable                            (mm_interconnect_0_nios2e_debug_mem_slave_byteenable),       //                                                       .byteenable
		.nios2e_debug_mem_slave_waitrequest                           (mm_interconnect_0_nios2e_debug_mem_slave_waitrequest),      //                                                       .waitrequest
		.nios2e_debug_mem_slave_debugaccess                           (mm_interconnect_0_nios2e_debug_mem_slave_debugaccess),      //                                                       .debugaccess
		.onchip_ram_s1_address                                        (mm_interconnect_0_onchip_ram_s1_address),                   //                                          onchip_ram_s1.address
		.onchip_ram_s1_write                                          (mm_interconnect_0_onchip_ram_s1_write),                     //                                                       .write
		.onchip_ram_s1_readdata                                       (mm_interconnect_0_onchip_ram_s1_readdata),                  //                                                       .readdata
		.onchip_ram_s1_writedata                                      (mm_interconnect_0_onchip_ram_s1_writedata),                 //                                                       .writedata
		.onchip_ram_s1_byteenable                                     (mm_interconnect_0_onchip_ram_s1_byteenable),                //                                                       .byteenable
		.onchip_ram_s1_chipselect                                     (mm_interconnect_0_onchip_ram_s1_chipselect),                //                                                       .chipselect
		.onchip_ram_s1_clken                                          (mm_interconnect_0_onchip_ram_s1_clken),                     //                                                       .clken
		.vga_out_slave_address                                        (mm_interconnect_0_vga_out_slave_address),                   //                                          vga_out_slave.address
		.vga_out_slave_write                                          (mm_interconnect_0_vga_out_slave_write),                     //                                                       .write
		.vga_out_slave_read                                           (mm_interconnect_0_vga_out_slave_read),                      //                                                       .read
		.vga_out_slave_readdata                                       (mm_interconnect_0_vga_out_slave_readdata),                  //                                                       .readdata
		.vga_out_slave_writedata                                      (mm_interconnect_0_vga_out_slave_writedata),                 //                                                       .writedata
		.vga_out_slave_waitrequest                                    (mm_interconnect_0_vga_out_slave_waitrequest)                //                                                       .waitrequest
	);

	pd_block_mm_interconnect_1 mm_interconnect_1 (
		.clock_clk_clk                                         (clock_clk),                                //                                       clock_clk.clk
		.bridge2_reset_reset_bridge_in_reset_reset             (rst_controller_reset_out_reset),           //             bridge2_reset_reset_bridge_in_reset.reset
		.frame_reader_clock_sreset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),           // frame_reader_clock_sreset_reset_bridge_in_reset.reset
		.bridge2_m0_address                                    (bridge2_m0_address),                       //                                      bridge2_m0.address
		.bridge2_m0_waitrequest                                (bridge2_m0_waitrequest),                   //                                                .waitrequest
		.bridge2_m0_burstcount                                 (bridge2_m0_burstcount),                    //                                                .burstcount
		.bridge2_m0_byteenable                                 (bridge2_m0_byteenable),                    //                                                .byteenable
		.bridge2_m0_read                                       (bridge2_m0_read),                          //                                                .read
		.bridge2_m0_readdata                                   (bridge2_m0_readdata),                      //                                                .readdata
		.bridge2_m0_readdatavalid                              (bridge2_m0_readdatavalid),                 //                                                .readdatavalid
		.bridge2_m0_write                                      (bridge2_m0_write),                         //                                                .write
		.bridge2_m0_writedata                                  (bridge2_m0_writedata),                     //                                                .writedata
		.bridge2_m0_debugaccess                                (bridge2_m0_debugaccess),                   //                                                .debugaccess
		.frame_reader_read_master_address                      (frame_reader_read_master_address),         //                        frame_reader_read_master.address
		.frame_reader_read_master_waitrequest                  (frame_reader_read_master_waitrequest),     //                                                .waitrequest
		.frame_reader_read_master_byteenable                   (frame_reader_read_master_byteenable),      //                                                .byteenable
		.frame_reader_read_master_read                         (frame_reader_read_master_read),            //                                                .read
		.frame_reader_read_master_readdata                     (frame_reader_read_master_readdata),        //                                                .readdata
		.frame_reader_read_master_readdatavalid                (frame_reader_read_master_readdatavalid),   //                                                .readdatavalid
		.sdram_s1_address                                      (mm_interconnect_1_sdram_s1_address),       //                                        sdram_s1.address
		.sdram_s1_write                                        (mm_interconnect_1_sdram_s1_write),         //                                                .write
		.sdram_s1_read                                         (mm_interconnect_1_sdram_s1_read),          //                                                .read
		.sdram_s1_readdata                                     (mm_interconnect_1_sdram_s1_readdata),      //                                                .readdata
		.sdram_s1_writedata                                    (mm_interconnect_1_sdram_s1_writedata),     //                                                .writedata
		.sdram_s1_byteenable                                   (mm_interconnect_1_sdram_s1_byteenable),    //                                                .byteenable
		.sdram_s1_readdatavalid                                (mm_interconnect_1_sdram_s1_readdatavalid), //                                                .readdatavalid
		.sdram_s1_waitrequest                                  (mm_interconnect_1_sdram_s1_waitrequest),   //                                                .waitrequest
		.sdram_s1_chipselect                                   (mm_interconnect_1_sdram_s1_chipselect)     //                                                .chipselect
	);

	pd_block_mm_interconnect_2 mm_interconnect_2 (
		.clock_clk_clk                                          (clock_clk),                                        //                                        clock_clk.clk
		.bridge1_reset_reset_bridge_in_reset_reset              (rst_controller_reset_out_reset),                   //              bridge1_reset_reset_bridge_in_reset.reset
		.dma_clock_sreset_reset_bridge_in_reset_reset           (rst_controller_002_reset_out_reset),               //           dma_clock_sreset_reset_bridge_in_reset.reset
		.dma_slave_translator_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),               // dma_slave_translator_reset_reset_bridge_in_reset.reset
		.rgb_tensor_reset_sink_reset_bridge_in_reset_reset      (rst_controller_reset_out_reset),                   //      rgb_tensor_reset_sink_reset_bridge_in_reset.reset
		.bridge1_m0_address                                     (bridge1_m0_address),                               //                                       bridge1_m0.address
		.bridge1_m0_waitrequest                                 (bridge1_m0_waitrequest),                           //                                                 .waitrequest
		.bridge1_m0_burstcount                                  (bridge1_m0_burstcount),                            //                                                 .burstcount
		.bridge1_m0_byteenable                                  (bridge1_m0_byteenable),                            //                                                 .byteenable
		.bridge1_m0_read                                        (bridge1_m0_read),                                  //                                                 .read
		.bridge1_m0_readdata                                    (bridge1_m0_readdata),                              //                                                 .readdata
		.bridge1_m0_readdatavalid                               (bridge1_m0_readdatavalid),                         //                                                 .readdatavalid
		.bridge1_m0_write                                       (bridge1_m0_write),                                 //                                                 .write
		.bridge1_m0_writedata                                   (bridge1_m0_writedata),                             //                                                 .writedata
		.bridge1_m0_debugaccess                                 (bridge1_m0_debugaccess),                           //                                                 .debugaccess
		.conv1_slave_address                                    (mm_interconnect_2_conv1_slave_address),            //                                      conv1_slave.address
		.conv1_slave_write                                      (mm_interconnect_2_conv1_slave_write),              //                                                 .write
		.conv1_slave_writedata                                  (mm_interconnect_2_conv1_slave_writedata),          //                                                 .writedata
		.conv1_slave_waitrequest                                (mm_interconnect_2_conv1_slave_waitrequest),        //                                                 .waitrequest
		.dma_slave_address                                      (mm_interconnect_2_dma_slave_address),              //                                        dma_slave.address
		.dma_slave_write                                        (mm_interconnect_2_dma_slave_write),                //                                                 .write
		.dma_slave_read                                         (mm_interconnect_2_dma_slave_read),                 //                                                 .read
		.dma_slave_readdata                                     (mm_interconnect_2_dma_slave_readdata),             //                                                 .readdata
		.dma_slave_writedata                                    (mm_interconnect_2_dma_slave_writedata),            //                                                 .writedata
		.dma_slave_waitrequest                                  (mm_interconnect_2_dma_slave_waitrequest),          //                                                 .waitrequest
		.from_memory1_slave_address                             (mm_interconnect_2_from_memory1_slave_address),     //                               from_memory1_slave.address
		.from_memory1_slave_write                               (mm_interconnect_2_from_memory1_slave_write),       //                                                 .write
		.from_memory1_slave_read                                (mm_interconnect_2_from_memory1_slave_read),        //                                                 .read
		.from_memory1_slave_readdata                            (mm_interconnect_2_from_memory1_slave_readdata),    //                                                 .readdata
		.from_memory1_slave_writedata                           (mm_interconnect_2_from_memory1_slave_writedata),   //                                                 .writedata
		.from_memory1_slave_waitrequest                         (mm_interconnect_2_from_memory1_slave_waitrequest), //                                                 .waitrequest
		.rgb_tensor_slave_address                               (mm_interconnect_2_rgb_tensor_slave_address),       //                                 rgb_tensor_slave.address
		.rgb_tensor_slave_write                                 (mm_interconnect_2_rgb_tensor_slave_write),         //                                                 .write
		.rgb_tensor_slave_read                                  (mm_interconnect_2_rgb_tensor_slave_read),          //                                                 .read
		.rgb_tensor_slave_readdata                              (mm_interconnect_2_rgb_tensor_slave_readdata),      //                                                 .readdata
		.rgb_tensor_slave_writedata                             (mm_interconnect_2_rgb_tensor_slave_writedata),     //                                                 .writedata
		.rgb_tensor_slave_waitrequest                           (mm_interconnect_2_rgb_tensor_slave_waitrequest)    //                                                 .waitrequest
	);

	pd_block_irq_mapper irq_mapper (
		.clk           (clock_clk),                      //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2e_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~clock_sreset_reset_n),              // reset_in0.reset
		.clk            (clock_clk),                          //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~clock_sreset_reset_n),              // reset_in0.reset
		.reset_in1      (nios2e_debug_reset_request_reset),   // reset_in1.reset
		.clk            (clock_clk),                          //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~clock_sreset_reset_n),              // reset_in0.reset
		.reset_in1      (nios2e_debug_reset_request_reset),   // reset_in1.reset
		.clk            (clock_clk),                          //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
