module sdram_input_efifo_module (
                                           // inputs:
                                            clock,
                                            rd,
                                            clock_sreset,
                                            wr,
                                            wr_data,

                                           // outputs:
                                            almost_empty,
                                            almost_full,
                                            empty,
                                            full,
                                            rd_data
                                         )
;

  output           almost_empty;
  output           almost_full;
  output           empty;
  output           full;
  output  [ 43: 0] rd_data;
  input            clock;
  input            rd;
  input            clock_sreset;
  input            wr;
  input   [ 43: 0] wr_data;


localparam ONE = 128'h1;
localparam ZERO = 128'h0;
  
wire             almost_empty;
wire             almost_full;
wire             empty;
reg     [  1: 0] entries;
reg     [ 43: 0] entry_0;
reg     [ 43: 0] entry_1;
wire             full;
reg              rd_address;
reg     [ 43: 0] rd_data;
wire    [  1: 0] rdwr;
reg              wr_address;
  assign rdwr = {rd, wr};
  assign full = entries == 2;
  assign almost_full = entries >= 1;
  assign empty = entries == 0;
  assign almost_empty = entries <= 1;
  always @(entry_0 or entry_1 or rd_address)
    begin
      case (rd_address) // synthesis parallel_case full_case
      
          1'd0: begin
              rd_data = entry_0;
          end // 1'd0 
      
          1'd1: begin
              rd_data = entry_1;
          end // 1'd1 
      
          //default: begin
          //end // default
      
      endcase // rd_address
    end


  always @(posedge clock)
    begin
      if (clock_sreset)
        begin
          wr_address <= 0;
          rd_address <= 0;
          entries <= 0;
        end
      else 
        case (rdwr) // synthesis parallel_case full_case
        
            2'd1: begin
                // Write data
                if (!full)
                  begin
                    entries <= entries + ONE[1:0];
                    wr_address <= (wr_address == ONE[0]) ? ZERO[0] : (wr_address + ONE[0]);
                  end
            end // 2'd1 
        
            2'd2: begin
                // Read data
                if (!empty)
                  begin
                    entries <= entries - ONE[1:0];
                    rd_address <= (rd_address == ONE[0]) ? ZERO[0] : (rd_address + ONE[1]);
                  end
            end // 2'd2 
        
            2'd3: begin
                wr_address <= (wr_address == 1) ? ZERO[0] : (wr_address + ONE[0]);
                rd_address <= (rd_address == 1) ? ZERO[0] : (rd_address + ONE[0]);
            end // 2'd3 
        
            //default: begin
            //end // default
        
        endcase // rdwr
    end


  always @(posedge clock)
    begin
      //Write data
      if (wr & !full)
          case (wr_address) // synthesis parallel_case full_case
          
              1'd0: begin
                  entry_0 <= wr_data;
              end // 1'd0 
          
              1'd1: begin
                  entry_1 <= wr_data;
              end // 1'd1 
          
              //default: begin
              //end // default
          
          endcase // wr_address
    end



endmodule
