// platform_designer_block.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module platform_designer_block (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire  [15:0] convolution_avalon_master_readdata;                        // mm_interconnect_0:convolution_avalon_master_readdata -> convolution:m_readdata
	wire         convolution_avalon_master_waitrequest;                     // mm_interconnect_0:convolution_avalon_master_waitrequest -> convolution:m_waitrequest
	wire  [31:0] convolution_avalon_master_address;                         // convolution:m_address -> mm_interconnect_0:convolution_avalon_master_address
	wire   [1:0] convolution_avalon_master_byteenable;                      // convolution:m_byteenable -> mm_interconnect_0:convolution_avalon_master_byteenable
	wire         convolution_avalon_master_read;                            // convolution:m_read -> mm_interconnect_0:convolution_avalon_master_read
	wire         convolution_avalon_master_readdatavalid;                   // mm_interconnect_0:convolution_avalon_master_readdatavalid -> convolution:m_readdatavalid
	wire  [15:0] convolution_avalon_master_writedata;                       // convolution:m_writedata -> mm_interconnect_0:convolution_avalon_master_writedata
	wire         convolution_avalon_master_write;                           // convolution:m_write -> mm_interconnect_0:convolution_avalon_master_write
	wire   [8:0] convolution_avalon_master_burstcount;                      // convolution:m_burstcount -> mm_interconnect_0:convolution_avalon_master_burstcount
	wire  [31:0] nios_data_master_readdata;                                 // mm_interconnect_0:nios_data_master_readdata -> nios:d_readdata
	wire         nios_data_master_waitrequest;                              // mm_interconnect_0:nios_data_master_waitrequest -> nios:d_waitrequest
	wire         nios_data_master_debugaccess;                              // nios:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios_data_master_debugaccess
	wire  [15:0] nios_data_master_address;                                  // nios:d_address -> mm_interconnect_0:nios_data_master_address
	wire   [3:0] nios_data_master_byteenable;                               // nios:d_byteenable -> mm_interconnect_0:nios_data_master_byteenable
	wire         nios_data_master_read;                                     // nios:d_read -> mm_interconnect_0:nios_data_master_read
	wire         nios_data_master_write;                                    // nios:d_write -> mm_interconnect_0:nios_data_master_write
	wire  [31:0] nios_data_master_writedata;                                // nios:d_writedata -> mm_interconnect_0:nios_data_master_writedata
	wire  [31:0] nios_instruction_master_readdata;                          // mm_interconnect_0:nios_instruction_master_readdata -> nios:i_readdata
	wire         nios_instruction_master_waitrequest;                       // mm_interconnect_0:nios_instruction_master_waitrequest -> nios:i_waitrequest
	wire  [15:0] nios_instruction_master_address;                           // nios:i_address -> mm_interconnect_0:nios_instruction_master_address
	wire         nios_instruction_master_read;                              // nios:i_read -> mm_interconnect_0:nios_instruction_master_read
	wire         mm_interconnect_0_onchip_ram_s1_chipselect;                // mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_readdata;                  // onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	wire  [12:0] mm_interconnect_0_onchip_ram_s1_address;                   // mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	wire   [3:0] mm_interconnect_0_onchip_ram_s1_byteenable;                // mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	wire         mm_interconnect_0_onchip_ram_s1_write;                     // mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_writedata;                 // mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	wire         mm_interconnect_0_onchip_ram_s1_clken;                     // mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_readdata;           // nios:debug_mem_slave_readdata -> mm_interconnect_0:nios_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_debug_mem_slave_waitrequest;        // nios:debug_mem_slave_waitrequest -> mm_interconnect_0:nios_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_debug_mem_slave_debugaccess;        // mm_interconnect_0:nios_debug_mem_slave_debugaccess -> nios:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_debug_mem_slave_address;            // mm_interconnect_0:nios_debug_mem_slave_address -> nios:debug_mem_slave_address
	wire         mm_interconnect_0_nios_debug_mem_slave_read;               // mm_interconnect_0:nios_debug_mem_slave_read -> nios:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_debug_mem_slave_byteenable;         // mm_interconnect_0:nios_debug_mem_slave_byteenable -> nios:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_debug_mem_slave_write;              // mm_interconnect_0:nios_debug_mem_slave_write -> nios:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_writedata;          // mm_interconnect_0:nios_debug_mem_slave_writedata -> nios:debug_mem_slave_writedata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_convolution_slave_readdata;              // convolution:s_readdata -> mm_interconnect_0:convolution_slave_readdata
	wire         mm_interconnect_0_convolution_slave_waitrequest;           // convolution:s_waitrequest -> mm_interconnect_0:convolution_slave_waitrequest
	wire   [3:0] mm_interconnect_0_convolution_slave_address;               // mm_interconnect_0:convolution_slave_address -> convolution:s_address
	wire         mm_interconnect_0_convolution_slave_read;                  // mm_interconnect_0:convolution_slave_read -> convolution:s_read
	wire         mm_interconnect_0_convolution_slave_write;                 // mm_interconnect_0:convolution_slave_write -> convolution:s_write
	wire  [31:0] mm_interconnect_0_convolution_slave_writedata;             // mm_interconnect_0:convolution_slave_writedata -> convolution:s_writedata
	wire         irq_mapper_receiver0_irq;                                  // convolution:s_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios_irq_irq;                                              // irq_mapper:sender_irq -> nios:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> convolution:clock_sreset
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:convolution_clock_sreset_reset_bridge_in_reset_reset, mm_interconnect_0:nios_reset_reset_bridge_in_reset_reset, nios:reset_n, onchip_ram:reset, rst_translator:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                    // rst_controller_001:reset_req -> [nios:reset_req, onchip_ram:reset_req, rst_translator:reset_req_in]

	convolution_burst #(
		.MAX_XRES    (34),
		.XRES1       (34),
		.XRES2       (18),
		.XRES3       (10),
		.XRES4       (6),
		.XRES5       (6),
		.YRES1       (34),
		.YRES2       (18),
		.YRES3       (10),
		.YRES4       (6),
		.YRES5       (6),
		.RESOLUTIONS (3),
		.KX          (3),
		.KY          (3),
		.EXP         (8),
		.MANT        (7),
		.WIDTHF      (16),
		.FIFO_DEPTH  (512),
		.WIDTH       (16),
		.WIDTHBE     (2),
		.WIDTHBC     (9)
	) convolution (
		.clock           (clk_clk),                                         //            clock.clk
		.clock_sreset    (rst_controller_reset_out_reset),                  //     clock_sreset.reset
		.s_address       (mm_interconnect_0_convolution_slave_address),     //            slave.address
		.s_writedata     (mm_interconnect_0_convolution_slave_writedata),   //                 .writedata
		.s_readdata      (mm_interconnect_0_convolution_slave_readdata),    //                 .readdata
		.s_read          (mm_interconnect_0_convolution_slave_read),        //                 .read
		.s_write         (mm_interconnect_0_convolution_slave_write),       //                 .write
		.s_waitrequest   (mm_interconnect_0_convolution_slave_waitrequest), //                 .waitrequest
		.m_address       (convolution_avalon_master_address),               //    avalon_master.address
		.m_readdata      (convolution_avalon_master_readdata),              //                 .readdata
		.m_writedata     (convolution_avalon_master_writedata),             //                 .writedata
		.m_byteenable    (convolution_avalon_master_byteenable),            //                 .byteenable
		.m_burstcount    (convolution_avalon_master_burstcount),            //                 .burstcount
		.m_read          (convolution_avalon_master_read),                  //                 .read
		.m_write         (convolution_avalon_master_write),                 //                 .write
		.m_readdatavalid (convolution_avalon_master_readdatavalid),         //                 .readdatavalid
		.m_waitrequest   (convolution_avalon_master_waitrequest),           //                 .waitrequest
		.s_irq           (irq_mapper_receiver0_irq)                         // interrupt_sender.irq
	);

	platform_designer_block_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	platform_designer_block_nios nios (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),             //                          .reset_req
		.d_address                           (nios_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_data_master_read),                              //                          .read
		.d_readdata                          (nios_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_data_master_write),                             //                          .write
		.d_writedata                         (nios_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                   //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	platform_designer_block_onchip_ram onchip_ram (
		.clk        (clk_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_onchip_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),     //       .reset_req
		.freeze     (1'b0)                                        // (terminated)
	);

	platform_designer_block_mm_interconnect_0 mm_interconnect_0 (
		.clock_clk_clk                                        (clk_clk),                                                   //                                      clock_clk.clk
		.convolution_clock_sreset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                        // convolution_clock_sreset_reset_bridge_in_reset.reset
		.nios_reset_reset_bridge_in_reset_reset               (rst_controller_001_reset_out_reset),                        //               nios_reset_reset_bridge_in_reset.reset
		.convolution_avalon_master_address                    (convolution_avalon_master_address),                         //                      convolution_avalon_master.address
		.convolution_avalon_master_waitrequest                (convolution_avalon_master_waitrequest),                     //                                               .waitrequest
		.convolution_avalon_master_burstcount                 (convolution_avalon_master_burstcount),                      //                                               .burstcount
		.convolution_avalon_master_byteenable                 (convolution_avalon_master_byteenable),                      //                                               .byteenable
		.convolution_avalon_master_read                       (convolution_avalon_master_read),                            //                                               .read
		.convolution_avalon_master_readdata                   (convolution_avalon_master_readdata),                        //                                               .readdata
		.convolution_avalon_master_readdatavalid              (convolution_avalon_master_readdatavalid),                   //                                               .readdatavalid
		.convolution_avalon_master_write                      (convolution_avalon_master_write),                           //                                               .write
		.convolution_avalon_master_writedata                  (convolution_avalon_master_writedata),                       //                                               .writedata
		.nios_data_master_address                             (nios_data_master_address),                                  //                               nios_data_master.address
		.nios_data_master_waitrequest                         (nios_data_master_waitrequest),                              //                                               .waitrequest
		.nios_data_master_byteenable                          (nios_data_master_byteenable),                               //                                               .byteenable
		.nios_data_master_read                                (nios_data_master_read),                                     //                                               .read
		.nios_data_master_readdata                            (nios_data_master_readdata),                                 //                                               .readdata
		.nios_data_master_write                               (nios_data_master_write),                                    //                                               .write
		.nios_data_master_writedata                           (nios_data_master_writedata),                                //                                               .writedata
		.nios_data_master_debugaccess                         (nios_data_master_debugaccess),                              //                                               .debugaccess
		.nios_instruction_master_address                      (nios_instruction_master_address),                           //                        nios_instruction_master.address
		.nios_instruction_master_waitrequest                  (nios_instruction_master_waitrequest),                       //                                               .waitrequest
		.nios_instruction_master_read                         (nios_instruction_master_read),                              //                                               .read
		.nios_instruction_master_readdata                     (nios_instruction_master_readdata),                          //                                               .readdata
		.convolution_slave_address                            (mm_interconnect_0_convolution_slave_address),               //                              convolution_slave.address
		.convolution_slave_write                              (mm_interconnect_0_convolution_slave_write),                 //                                               .write
		.convolution_slave_read                               (mm_interconnect_0_convolution_slave_read),                  //                                               .read
		.convolution_slave_readdata                           (mm_interconnect_0_convolution_slave_readdata),              //                                               .readdata
		.convolution_slave_writedata                          (mm_interconnect_0_convolution_slave_writedata),             //                                               .writedata
		.convolution_slave_waitrequest                        (mm_interconnect_0_convolution_slave_waitrequest),           //                                               .waitrequest
		.jtag_uart_avalon_jtag_slave_address                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                    jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                               .write
		.jtag_uart_avalon_jtag_slave_read                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                               .read
		.jtag_uart_avalon_jtag_slave_readdata                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                               .readdata
		.jtag_uart_avalon_jtag_slave_writedata                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                               .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                               .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                               .chipselect
		.nios_debug_mem_slave_address                         (mm_interconnect_0_nios_debug_mem_slave_address),            //                           nios_debug_mem_slave.address
		.nios_debug_mem_slave_write                           (mm_interconnect_0_nios_debug_mem_slave_write),              //                                               .write
		.nios_debug_mem_slave_read                            (mm_interconnect_0_nios_debug_mem_slave_read),               //                                               .read
		.nios_debug_mem_slave_readdata                        (mm_interconnect_0_nios_debug_mem_slave_readdata),           //                                               .readdata
		.nios_debug_mem_slave_writedata                       (mm_interconnect_0_nios_debug_mem_slave_writedata),          //                                               .writedata
		.nios_debug_mem_slave_byteenable                      (mm_interconnect_0_nios_debug_mem_slave_byteenable),         //                                               .byteenable
		.nios_debug_mem_slave_waitrequest                     (mm_interconnect_0_nios_debug_mem_slave_waitrequest),        //                                               .waitrequest
		.nios_debug_mem_slave_debugaccess                     (mm_interconnect_0_nios_debug_mem_slave_debugaccess),        //                                               .debugaccess
		.onchip_ram_s1_address                                (mm_interconnect_0_onchip_ram_s1_address),                   //                                  onchip_ram_s1.address
		.onchip_ram_s1_write                                  (mm_interconnect_0_onchip_ram_s1_write),                     //                                               .write
		.onchip_ram_s1_readdata                               (mm_interconnect_0_onchip_ram_s1_readdata),                  //                                               .readdata
		.onchip_ram_s1_writedata                              (mm_interconnect_0_onchip_ram_s1_writedata),                 //                                               .writedata
		.onchip_ram_s1_byteenable                             (mm_interconnect_0_onchip_ram_s1_byteenable),                //                                               .byteenable
		.onchip_ram_s1_chipselect                             (mm_interconnect_0_onchip_ram_s1_chipselect),                //                                               .chipselect
		.onchip_ram_s1_clken                                  (mm_interconnect_0_onchip_ram_s1_clken)                      //                                               .clken
	);

	platform_designer_block_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (nios_irq_irq)                        //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
