// internal_oscillator.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module internal_oscillator (
		output wire  clkout, // clkout.clk
		input  wire  oscena  // oscena.oscena
	);

	altera_int_osc int_osc_0 (
		.oscena (oscena), // oscena.oscena
		.clkout (clkout)  // clkout.clk
	);

endmodule
