
module internal_oscillator (
	clkout,
	oscena);	

	output		clkout;
	input		oscena;
endmodule
