
module internal_oscillator (
	oscena,
	clkout);	

	input		oscena;
	output		clkout;
endmodule
