// recursive module function powers of two only (for now)
module fp_add_tree # (
            parameter                       EXP = 8,
            parameter                       MANT = 7,
            parameter                       ITEMS = 32,
            parameter                       WIDTH = 1 + EXP + MANT,
            parameter                       EXTRA_PIPELINE = 0
)
(
    input   logic                           clock,
    input   logic                           clock_sreset,
    input   logic                           data_valid,
    input   logic [ITEMS-1:0][WIDTH-1:0]    data,
    output  logic                           result_valid,
    output  logic [WIDTH-1:0]               result
);
            localparam                      HALF = (ITEMS / 2);
            localparam                      WIDTHH = (ITEMS - HALF);
            localparam                      ZERO = {WIDTH{1'b0}};
    generate
        begin
            if (ITEMS == 2) begin   // only one branch?
                fp_add                     # (
                                                .EXP(EXP),
                                                .MANT(MANT),
                                                .WIDTH(WIDTH),
                                                .EXTRA_PIPELINE(EXTRA_PIPELINE)
                                            )
                                            addera (
                                                .clock(clock),
                                                .clock_sreset(clock_sreset),
                                                .data_valid(data_valid),
                                                .dataa(data[0]),
                                                .datab(data[1]),
                                                .result_valid(result_valid),
                                                .result(result)
                                            );
            end
            if (ITEMS > 2) begin // keep halving the tree
                logic [WIDTH-1:0]           resulta, resultb;
                logic                       resulta_valid;
                fp_add_tree                 # (
                                                .EXP(EXP),
                                                .MANT(MANT),
                                                .ITEMS(HALF),
                                                .EXTRA_PIPELINE(EXTRA_PIPELINE)
                                            )
                                            addera (
                                                .clock(clock),
                                                .clock_sreset(clock_sreset),
                                                .data_valid(data_valid),
                                                .data(data[ITEMS-1:WIDTHH]),
                                                .result_valid(resulta_valid),
                                                .result(resulta)
                                            );
                fp_add_tree                 # (
                                                .EXP(EXP),
                                                .MANT(MANT),
                                                .ITEMS(WIDTHH),
                                                .EXTRA_PIPELINE(EXTRA_PIPELINE)
                                            )
                                            adderb (
                                                .clock(clock),
                                                .clock_sreset(clock_sreset),
                                                .data_valid(),
                                                .data(data[WIDTHH-1:0]),
                                                .result_valid(),
                                                .result(resultb)
                                            );
                fp_add                      # (
                                                .EXP(EXP),
                                                .MANT(MANT),
                                                .WIDTH(WIDTH),
                                                .EXTRA_PIPELINE(EXTRA_PIPELINE)
                                            )
                                            adderc (
                                                .clock(clock),
                                                .clock_sreset(clock_sreset),
                                                .data_valid(resulta_valid),
                                                .dataa(resulta),
                                                .datab(resultb),
                                                .result_valid(result_valid),
                                                .result(result)
                                            );
         end
      end
   endgenerate

endmodule
