// pd_block.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module pd_block (
		input  wire        clock_clk,                //            clock.clk
		input  wire        clock_sreset_reset_n,     //     clock_sreset.reset_n
		output wire [9:0]  led_export,               //              led.export
		output wire [12:0] sdram_addr,               //            sdram.addr
		output wire [1:0]  sdram_ba,                 //                 .ba
		output wire        sdram_cas_n,              //                 .cas_n
		output wire        sdram_cke,                //                 .cke
		output wire        sdram_cs_n,               //                 .cs_n
		inout  wire [15:0] sdram_dq,                 //                 .dq
		output wire [1:0]  sdram_dqm,                //                 .dqm
		output wire        sdram_ras_n,              //                 .ras_n
		output wire        sdram_we_n,               //                 .we_n
		input  wire        vga_clock_clk,            //        vga_clock.clk
		input  wire        vga_clock_sreset_reset_n  // vga_clock_sreset.reset_n
	);

	wire  [15:0] convolution0_avalon_master_readdata;                       // mm_interconnect_0:convolution0_avalon_master_readdata -> convolution0:m_readdata
	wire         convolution0_avalon_master_waitrequest;                    // mm_interconnect_0:convolution0_avalon_master_waitrequest -> convolution0:m_waitrequest
	wire  [31:0] convolution0_avalon_master_address;                        // convolution0:m_address -> mm_interconnect_0:convolution0_avalon_master_address
	wire   [1:0] convolution0_avalon_master_byteenable;                     // convolution0:m_byteenable -> mm_interconnect_0:convolution0_avalon_master_byteenable
	wire         convolution0_avalon_master_read;                           // convolution0:m_read -> mm_interconnect_0:convolution0_avalon_master_read
	wire         convolution0_avalon_master_readdatavalid;                  // mm_interconnect_0:convolution0_avalon_master_readdatavalid -> convolution0:m_readdatavalid
	wire  [15:0] convolution0_avalon_master_writedata;                      // convolution0:m_writedata -> mm_interconnect_0:convolution0_avalon_master_writedata
	wire         convolution0_avalon_master_write;                          // convolution0:m_write -> mm_interconnect_0:convolution0_avalon_master_write
	wire   [8:0] convolution0_avalon_master_burstcount;                     // convolution0:m_burstcount -> mm_interconnect_0:convolution0_avalon_master_burstcount
	wire  [15:0] rgb_to_tensor_avalon_master_readdata;                      // mm_interconnect_0:rgb_to_tensor_avalon_master_readdata -> rgb_to_tensor:m_readdata
	wire         rgb_to_tensor_avalon_master_waitrequest;                   // mm_interconnect_0:rgb_to_tensor_avalon_master_waitrequest -> rgb_to_tensor:m_waitrequest
	wire  [31:0] rgb_to_tensor_avalon_master_address;                       // rgb_to_tensor:m_address -> mm_interconnect_0:rgb_to_tensor_avalon_master_address
	wire   [1:0] rgb_to_tensor_avalon_master_byteenable;                    // rgb_to_tensor:m_byteenable -> mm_interconnect_0:rgb_to_tensor_avalon_master_byteenable
	wire         rgb_to_tensor_avalon_master_read;                          // rgb_to_tensor:m_read -> mm_interconnect_0:rgb_to_tensor_avalon_master_read
	wire  [15:0] rgb_to_tensor_avalon_master_writedata;                     // rgb_to_tensor:m_writedata -> mm_interconnect_0:rgb_to_tensor_avalon_master_writedata
	wire         rgb_to_tensor_avalon_master_write;                         // rgb_to_tensor:m_write -> mm_interconnect_0:rgb_to_tensor_avalon_master_write
	wire  [31:0] nios2e_data_master_readdata;                               // mm_interconnect_0:nios2e_data_master_readdata -> nios2e:d_readdata
	wire         nios2e_data_master_waitrequest;                            // mm_interconnect_0:nios2e_data_master_waitrequest -> nios2e:d_waitrequest
	wire         nios2e_data_master_debugaccess;                            // nios2e:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2e_data_master_debugaccess
	wire  [26:0] nios2e_data_master_address;                                // nios2e:d_address -> mm_interconnect_0:nios2e_data_master_address
	wire   [3:0] nios2e_data_master_byteenable;                             // nios2e:d_byteenable -> mm_interconnect_0:nios2e_data_master_byteenable
	wire         nios2e_data_master_read;                                   // nios2e:d_read -> mm_interconnect_0:nios2e_data_master_read
	wire         nios2e_data_master_write;                                  // nios2e:d_write -> mm_interconnect_0:nios2e_data_master_write
	wire  [31:0] nios2e_data_master_writedata;                              // nios2e:d_writedata -> mm_interconnect_0:nios2e_data_master_writedata
	wire  [31:0] nios2e_instruction_master_readdata;                        // mm_interconnect_0:nios2e_instruction_master_readdata -> nios2e:i_readdata
	wire         nios2e_instruction_master_waitrequest;                     // mm_interconnect_0:nios2e_instruction_master_waitrequest -> nios2e:i_waitrequest
	wire  [26:0] nios2e_instruction_master_address;                         // nios2e:i_address -> mm_interconnect_0:nios2e_instruction_master_address
	wire         nios2e_instruction_master_read;                            // nios2e:i_read -> mm_interconnect_0:nios2e_instruction_master_read
	wire         mm_interconnect_0_sdram_s1_chipselect;                     // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                       // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                    // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                        // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                           // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                     // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                  // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                          // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                      // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [31:0] mm_interconnect_0_nios2e_debug_mem_slave_readdata;         // nios2e:debug_mem_slave_readdata -> mm_interconnect_0:nios2e_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2e_debug_mem_slave_waitrequest;      // nios2e:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2e_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2e_debug_mem_slave_debugaccess;      // mm_interconnect_0:nios2e_debug_mem_slave_debugaccess -> nios2e:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2e_debug_mem_slave_address;          // mm_interconnect_0:nios2e_debug_mem_slave_address -> nios2e:debug_mem_slave_address
	wire         mm_interconnect_0_nios2e_debug_mem_slave_read;             // mm_interconnect_0:nios2e_debug_mem_slave_read -> nios2e:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2e_debug_mem_slave_byteenable;       // mm_interconnect_0:nios2e_debug_mem_slave_byteenable -> nios2e:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2e_debug_mem_slave_write;            // mm_interconnect_0:nios2e_debug_mem_slave_write -> nios2e:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2e_debug_mem_slave_writedata;        // mm_interconnect_0:nios2e_debug_mem_slave_writedata -> nios2e:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_ram_s1_chipselect;                // mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_readdata;                  // onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	wire  [11:0] mm_interconnect_0_onchip_ram_s1_address;                   // mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	wire   [3:0] mm_interconnect_0_onchip_ram_s1_byteenable;                // mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	wire         mm_interconnect_0_onchip_ram_s1_write;                     // mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_writedata;                 // mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	wire         mm_interconnect_0_onchip_ram_s1_clken;                     // mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_convolution0_avalon_slave_readdata;      // convolution0:s_readdata -> mm_interconnect_0:convolution0_avalon_slave_readdata
	wire         mm_interconnect_0_convolution0_avalon_slave_waitrequest;   // convolution0:s_waitrequest -> mm_interconnect_0:convolution0_avalon_slave_waitrequest
	wire   [3:0] mm_interconnect_0_convolution0_avalon_slave_address;       // mm_interconnect_0:convolution0_avalon_slave_address -> convolution0:s_address
	wire         mm_interconnect_0_convolution0_avalon_slave_read;          // mm_interconnect_0:convolution0_avalon_slave_read -> convolution0:s_read
	wire         mm_interconnect_0_convolution0_avalon_slave_write;         // mm_interconnect_0:convolution0_avalon_slave_write -> convolution0:s_write
	wire  [31:0] mm_interconnect_0_convolution0_avalon_slave_writedata;     // mm_interconnect_0:convolution0_avalon_slave_writedata -> convolution0:s_writedata
	wire         mm_interconnect_0_led_s1_chipselect;                       // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                         // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;                          // mm_interconnect_0:led_s1_address -> led:address
	wire         mm_interconnect_0_led_s1_write;                            // mm_interconnect_0:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                        // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire  [31:0] mm_interconnect_0_rgb_to_tensor_slave_readdata;            // rgb_to_tensor:s_readdata -> mm_interconnect_0:rgb_to_tensor_slave_readdata
	wire         mm_interconnect_0_rgb_to_tensor_slave_waitrequest;         // rgb_to_tensor:s_waitrequest -> mm_interconnect_0:rgb_to_tensor_slave_waitrequest
	wire   [3:0] mm_interconnect_0_rgb_to_tensor_slave_address;             // mm_interconnect_0:rgb_to_tensor_slave_address -> rgb_to_tensor:s_address
	wire         mm_interconnect_0_rgb_to_tensor_slave_read;                // mm_interconnect_0:rgb_to_tensor_slave_read -> rgb_to_tensor:s_read
	wire         mm_interconnect_0_rgb_to_tensor_slave_write;               // mm_interconnect_0:rgb_to_tensor_slave_write -> rgb_to_tensor:s_write
	wire  [31:0] mm_interconnect_0_rgb_to_tensor_slave_writedata;           // mm_interconnect_0:rgb_to_tensor_slave_writedata -> rgb_to_tensor:s_writedata
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2e_irq_irq;                                            // irq_mapper:sender_irq -> nios2e:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [irq_mapper:reset, jtag_uart:rst_n, led:reset_n, mm_interconnect_0:convolution0_clock_sreset_reset_bridge_in_reset_reset, mm_interconnect_0:nios2e_reset_reset_bridge_in_reset_reset, nios2e:reset_n, onchip_ram:reset, rst_translator:in_reset, sdram:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [nios2e:reset_req, onchip_ram:reset_req, rst_translator:reset_req_in]

	convolution_burst #(
		.MAX_RES        (256),
		.XRES1          (16),
		.XRES2          (32),
		.XRES3          (64),
		.XRES4          (128),
		.XRES5          (256),
		.YRES1          (16),
		.YRES2          (32),
		.YRES3          (64),
		.YRES4          (128),
		.YRES5          (256),
		.RESOLUTIONS    (5),
		.PAD            (1),
		.KX             (3),
		.KY             (3),
		.EXP            (8),
		.MANT           (7),
		.WIDTHF         (16),
		.FIFO_DEPTH     (512),
		.WIDTH          (16),
		.WIDTHB         (2),
		.WIDTHD         (9),
		.ADDER_PIPELINE (1)
	) convolution0 (
		.m_address       (convolution0_avalon_master_address),                      // avalon_master.address
		.m_readdata      (convolution0_avalon_master_readdata),                     //              .readdata
		.m_writedata     (convolution0_avalon_master_writedata),                    //              .writedata
		.m_byteenable    (convolution0_avalon_master_byteenable),                   //              .byteenable
		.m_burstcount    (convolution0_avalon_master_burstcount),                   //              .burstcount
		.m_read          (convolution0_avalon_master_read),                         //              .read
		.m_write         (convolution0_avalon_master_write),                        //              .write
		.m_readdatavalid (convolution0_avalon_master_readdatavalid),                //              .readdatavalid
		.m_waitrequest   (convolution0_avalon_master_waitrequest),                  //              .waitrequest
		.s_address       (mm_interconnect_0_convolution0_avalon_slave_address),     //  avalon_slave.address
		.s_writedata     (mm_interconnect_0_convolution0_avalon_slave_writedata),   //              .writedata
		.s_readdata      (mm_interconnect_0_convolution0_avalon_slave_readdata),    //              .readdata
		.s_read          (mm_interconnect_0_convolution0_avalon_slave_read),        //              .read
		.s_write         (mm_interconnect_0_convolution0_avalon_slave_write),       //              .write
		.s_waitrequest   (mm_interconnect_0_convolution0_avalon_slave_waitrequest), //              .waitrequest
		.clock           (clock_clk),                                               //         clock.clk
		.clock_sreset    (~clock_sreset_reset_n)                                    //  clock_sreset.reset
	);

	pd_block_jtag_uart jtag_uart (
		.clk            (clock_clk),                                                 //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	pd_block_led led (
		.clk        (clock_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                           // external_connection.export
	);

	pd_block_nios2e nios2e (
		.clk                                 (clock_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (nios2e_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2e_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2e_data_master_read),                              //                          .read
		.d_readdata                          (nios2e_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2e_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2e_data_master_write),                             //                          .write
		.d_writedata                         (nios2e_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2e_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2e_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2e_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2e_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2e_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2e_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2e_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2e_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2e_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2e_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2e_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2e_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2e_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2e_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                      // custom_instruction_master.readra
	);

	pd_block_onchip_ram onchip_ram (
		.clk        (clock_clk),                                  //   clk1.clk
		.address    (mm_interconnect_0_onchip_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                        // (terminated)
	);

	rgb_to_tensor rgb_to_tensor (
		.s_address     (mm_interconnect_0_rgb_to_tensor_slave_address),     //         slave.address
		.s_readdata    (mm_interconnect_0_rgb_to_tensor_slave_readdata),    //              .readdata
		.s_writedata   (mm_interconnect_0_rgb_to_tensor_slave_writedata),   //              .writedata
		.s_read        (mm_interconnect_0_rgb_to_tensor_slave_read),        //              .read
		.s_write       (mm_interconnect_0_rgb_to_tensor_slave_write),       //              .write
		.s_waitrequest (mm_interconnect_0_rgb_to_tensor_slave_waitrequest), //              .waitrequest
		.m_address     (rgb_to_tensor_avalon_master_address),               // avalon_master.address
		.m_writedata   (rgb_to_tensor_avalon_master_writedata),             //              .writedata
		.m_readdata    (rgb_to_tensor_avalon_master_readdata),              //              .readdata
		.m_byteenable  (rgb_to_tensor_avalon_master_byteenable),            //              .byteenable
		.m_read        (rgb_to_tensor_avalon_master_read),                  //              .read
		.m_write       (rgb_to_tensor_avalon_master_write),                 //              .write
		.m_waitrequest (rgb_to_tensor_avalon_master_waitrequest),           //              .waitrequest
		.clock         (clock_clk),                                         //    clock_sink.clk
		.clock_sreset  (~clock_sreset_reset_n)                              //    reset_sink.reset
	);

	pd_block_sdram sdram (
		.clk            (clock_clk),                                //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	pd_block_mm_interconnect_0 mm_interconnect_0 (
		.clock_clk_clk                                         (clock_clk),                                                 //                                       clock_clk.clk
		.convolution0_clock_sreset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // convolution0_clock_sreset_reset_bridge_in_reset.reset
		.nios2e_reset_reset_bridge_in_reset_reset              (rst_controller_reset_out_reset),                            //              nios2e_reset_reset_bridge_in_reset.reset
		.convolution0_avalon_master_address                    (convolution0_avalon_master_address),                        //                      convolution0_avalon_master.address
		.convolution0_avalon_master_waitrequest                (convolution0_avalon_master_waitrequest),                    //                                                .waitrequest
		.convolution0_avalon_master_burstcount                 (convolution0_avalon_master_burstcount),                     //                                                .burstcount
		.convolution0_avalon_master_byteenable                 (convolution0_avalon_master_byteenable),                     //                                                .byteenable
		.convolution0_avalon_master_read                       (convolution0_avalon_master_read),                           //                                                .read
		.convolution0_avalon_master_readdata                   (convolution0_avalon_master_readdata),                       //                                                .readdata
		.convolution0_avalon_master_readdatavalid              (convolution0_avalon_master_readdatavalid),                  //                                                .readdatavalid
		.convolution0_avalon_master_write                      (convolution0_avalon_master_write),                          //                                                .write
		.convolution0_avalon_master_writedata                  (convolution0_avalon_master_writedata),                      //                                                .writedata
		.nios2e_data_master_address                            (nios2e_data_master_address),                                //                              nios2e_data_master.address
		.nios2e_data_master_waitrequest                        (nios2e_data_master_waitrequest),                            //                                                .waitrequest
		.nios2e_data_master_byteenable                         (nios2e_data_master_byteenable),                             //                                                .byteenable
		.nios2e_data_master_read                               (nios2e_data_master_read),                                   //                                                .read
		.nios2e_data_master_readdata                           (nios2e_data_master_readdata),                               //                                                .readdata
		.nios2e_data_master_write                              (nios2e_data_master_write),                                  //                                                .write
		.nios2e_data_master_writedata                          (nios2e_data_master_writedata),                              //                                                .writedata
		.nios2e_data_master_debugaccess                        (nios2e_data_master_debugaccess),                            //                                                .debugaccess
		.nios2e_instruction_master_address                     (nios2e_instruction_master_address),                         //                       nios2e_instruction_master.address
		.nios2e_instruction_master_waitrequest                 (nios2e_instruction_master_waitrequest),                     //                                                .waitrequest
		.nios2e_instruction_master_read                        (nios2e_instruction_master_read),                            //                                                .read
		.nios2e_instruction_master_readdata                    (nios2e_instruction_master_readdata),                        //                                                .readdata
		.rgb_to_tensor_avalon_master_address                   (rgb_to_tensor_avalon_master_address),                       //                     rgb_to_tensor_avalon_master.address
		.rgb_to_tensor_avalon_master_waitrequest               (rgb_to_tensor_avalon_master_waitrequest),                   //                                                .waitrequest
		.rgb_to_tensor_avalon_master_byteenable                (rgb_to_tensor_avalon_master_byteenable),                    //                                                .byteenable
		.rgb_to_tensor_avalon_master_read                      (rgb_to_tensor_avalon_master_read),                          //                                                .read
		.rgb_to_tensor_avalon_master_readdata                  (rgb_to_tensor_avalon_master_readdata),                      //                                                .readdata
		.rgb_to_tensor_avalon_master_write                     (rgb_to_tensor_avalon_master_write),                         //                                                .write
		.rgb_to_tensor_avalon_master_writedata                 (rgb_to_tensor_avalon_master_writedata),                     //                                                .writedata
		.convolution0_avalon_slave_address                     (mm_interconnect_0_convolution0_avalon_slave_address),       //                       convolution0_avalon_slave.address
		.convolution0_avalon_slave_write                       (mm_interconnect_0_convolution0_avalon_slave_write),         //                                                .write
		.convolution0_avalon_slave_read                        (mm_interconnect_0_convolution0_avalon_slave_read),          //                                                .read
		.convolution0_avalon_slave_readdata                    (mm_interconnect_0_convolution0_avalon_slave_readdata),      //                                                .readdata
		.convolution0_avalon_slave_writedata                   (mm_interconnect_0_convolution0_avalon_slave_writedata),     //                                                .writedata
		.convolution0_avalon_slave_waitrequest                 (mm_interconnect_0_convolution0_avalon_slave_waitrequest),   //                                                .waitrequest
		.jtag_uart_avalon_jtag_slave_address                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                                .write
		.jtag_uart_avalon_jtag_slave_read                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                                .read
		.jtag_uart_avalon_jtag_slave_readdata                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                                .chipselect
		.led_s1_address                                        (mm_interconnect_0_led_s1_address),                          //                                          led_s1.address
		.led_s1_write                                          (mm_interconnect_0_led_s1_write),                            //                                                .write
		.led_s1_readdata                                       (mm_interconnect_0_led_s1_readdata),                         //                                                .readdata
		.led_s1_writedata                                      (mm_interconnect_0_led_s1_writedata),                        //                                                .writedata
		.led_s1_chipselect                                     (mm_interconnect_0_led_s1_chipselect),                       //                                                .chipselect
		.nios2e_debug_mem_slave_address                        (mm_interconnect_0_nios2e_debug_mem_slave_address),          //                          nios2e_debug_mem_slave.address
		.nios2e_debug_mem_slave_write                          (mm_interconnect_0_nios2e_debug_mem_slave_write),            //                                                .write
		.nios2e_debug_mem_slave_read                           (mm_interconnect_0_nios2e_debug_mem_slave_read),             //                                                .read
		.nios2e_debug_mem_slave_readdata                       (mm_interconnect_0_nios2e_debug_mem_slave_readdata),         //                                                .readdata
		.nios2e_debug_mem_slave_writedata                      (mm_interconnect_0_nios2e_debug_mem_slave_writedata),        //                                                .writedata
		.nios2e_debug_mem_slave_byteenable                     (mm_interconnect_0_nios2e_debug_mem_slave_byteenable),       //                                                .byteenable
		.nios2e_debug_mem_slave_waitrequest                    (mm_interconnect_0_nios2e_debug_mem_slave_waitrequest),      //                                                .waitrequest
		.nios2e_debug_mem_slave_debugaccess                    (mm_interconnect_0_nios2e_debug_mem_slave_debugaccess),      //                                                .debugaccess
		.onchip_ram_s1_address                                 (mm_interconnect_0_onchip_ram_s1_address),                   //                                   onchip_ram_s1.address
		.onchip_ram_s1_write                                   (mm_interconnect_0_onchip_ram_s1_write),                     //                                                .write
		.onchip_ram_s1_readdata                                (mm_interconnect_0_onchip_ram_s1_readdata),                  //                                                .readdata
		.onchip_ram_s1_writedata                               (mm_interconnect_0_onchip_ram_s1_writedata),                 //                                                .writedata
		.onchip_ram_s1_byteenable                              (mm_interconnect_0_onchip_ram_s1_byteenable),                //                                                .byteenable
		.onchip_ram_s1_chipselect                              (mm_interconnect_0_onchip_ram_s1_chipselect),                //                                                .chipselect
		.onchip_ram_s1_clken                                   (mm_interconnect_0_onchip_ram_s1_clken),                     //                                                .clken
		.rgb_to_tensor_slave_address                           (mm_interconnect_0_rgb_to_tensor_slave_address),             //                             rgb_to_tensor_slave.address
		.rgb_to_tensor_slave_write                             (mm_interconnect_0_rgb_to_tensor_slave_write),               //                                                .write
		.rgb_to_tensor_slave_read                              (mm_interconnect_0_rgb_to_tensor_slave_read),                //                                                .read
		.rgb_to_tensor_slave_readdata                          (mm_interconnect_0_rgb_to_tensor_slave_readdata),            //                                                .readdata
		.rgb_to_tensor_slave_writedata                         (mm_interconnect_0_rgb_to_tensor_slave_writedata),           //                                                .writedata
		.rgb_to_tensor_slave_waitrequest                       (mm_interconnect_0_rgb_to_tensor_slave_waitrequest),         //                                                .waitrequest
		.sdram_s1_address                                      (mm_interconnect_0_sdram_s1_address),                        //                                        sdram_s1.address
		.sdram_s1_write                                        (mm_interconnect_0_sdram_s1_write),                          //                                                .write
		.sdram_s1_read                                         (mm_interconnect_0_sdram_s1_read),                           //                                                .read
		.sdram_s1_readdata                                     (mm_interconnect_0_sdram_s1_readdata),                       //                                                .readdata
		.sdram_s1_writedata                                    (mm_interconnect_0_sdram_s1_writedata),                      //                                                .writedata
		.sdram_s1_byteenable                                   (mm_interconnect_0_sdram_s1_byteenable),                     //                                                .byteenable
		.sdram_s1_readdatavalid                                (mm_interconnect_0_sdram_s1_readdatavalid),                  //                                                .readdatavalid
		.sdram_s1_waitrequest                                  (mm_interconnect_0_sdram_s1_waitrequest),                    //                                                .waitrequest
		.sdram_s1_chipselect                                   (mm_interconnect_0_sdram_s1_chipselect)                      //                                                .chipselect
	);

	pd_block_irq_mapper irq_mapper (
		.clk           (clock_clk),                      //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2e_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~clock_sreset_reset_n),              // reset_in0.reset
		.clk            (clock_clk),                          //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
