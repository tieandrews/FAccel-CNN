module bcd_mult16 (
    input   logic               clock,
    input   logic [15:0]        dataa,
    input   logic [15:0]        datab,
    output  logic [31:0]        result
);

    

endmodule
