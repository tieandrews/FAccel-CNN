
module oscillator (
	clkout,
	oscena);	

	output		clkout;
	input		oscena;
endmodule
